// Code your design he
	



      



